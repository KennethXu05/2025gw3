module wave_top#(
  parameter H_Visible_area    = 800, //��Ļ��ʾ������
  parameter V_Visible_area    = 480, //��Ļ��ʾ����߶�
  parameter H2_ActiveSize  =   750,
  parameter V2_ActiveSize  =   256
)(
  input clk,
  input clk_ctrl,
  input reset_n,
  //char_disp_hbegin,
  //char_disp_vbegin,
  input Frame_Begin,
  input [11:0]visible_hcount,
  input [11:0]visible_vcount,
  //ƫ������ԭ�㣨���Ͻǣ�  
  input  [11:0]   I_vtc2_offset_x,//�����Ļԭ��(���Ͻ�)X����ƫ��
  input  [11:0]   I_vtc2_offset_y,//�����Ļԭ��(���Ͻ�)Y����ƫ��
  //ͨ��1
  input I_wave1_clk,//����ʱ��1
  input [7:0] I_wave1_data,//��������1
  input I_wave1_data_de,//����������Ч1
  //ͨ��2
  input I_wave2_clk,//����ʱ��2
  input [7:0] I_wave2_data,//��������2
  input I_wave2_data_de,//����������Ч2

  input I_vtc_vs,
  input I_vtc_hs,
  input I_vtc_de,

  output reg O_vtc_vs,
  output reg O_vtc_hs,
  output reg O_vtc_de,
  output [15:0]O_vtc_rgb,

  input  single,
  
  input trigger_edge,//switch
  input trigger_button//button
  
);
    wire trigger_button_minus_flag;
    key_filter_wave key_filter_wave_single(
	.clk(clk),
	.reset_n(reset_n),

	.key_in(single),
	.key_flag(),
	.key_state(key_state)
);
    key_filter_wave key_filter_wave_trigger_button(
	.clk(clk),
	.reset_n(reset_n),

	.key_in(trigger_button),
	.key_flag(trigger_button_minus_flag),
	.key_state(trigger_button_state)
);
    key_filter_wave key_filter_wave_trigger_edge(
	.clk(clk),
	.reset_n(reset_n),

	.key_in(trigger_edge),
	.key_flag(),
	.key_state(trigger_edge_state)
);
    reg r_key_state;
    always @(posedge clk or negedge reset_n) begin
        if(!reset_n)
            r_key_state<=1;
        else
            r_key_state<=key_state;
    end
    reg single_flag;
    always @(posedge clk or negedge reset_n) begin
        if(!reset_n)
            single_flag<=0;
        else if({r_key_state,key_state}==2'b10)
            single_flag<=!single_flag;
        else
            single_flag<=single_flag;
    end
//trigger_button
    reg r_trigger_button_state;
    always @(posedge clk or negedge reset_n) begin
        if(!reset_n)
            r_trigger_button_state<=1;
        else
            r_trigger_button_state<=trigger_button_state;
    end
    reg trigger_button_flag;
    always @(posedge clk or negedge reset_n) begin
        if(!reset_n)
            trigger_button_flag<=0;
        else if({r_trigger_button_state,trigger_button_state}==2'b10)
            trigger_button_flag<=!trigger_button_flag;
        else
            trigger_button_flag<=trigger_button_flag;
    end
    //trigger_edge
        reg r_trigger_edge_state;
    always @(posedge clk or negedge reset_n) begin
        if(!reset_n)
            r_trigger_edge_state<=1;
        else
            r_trigger_edge_state<=trigger_edge_state;
    end
    reg trigger_edge_o;
    always @(posedge clk or negedge reset_n) begin
        if(!reset_n)
            trigger_edge_o<=0;
        else if({r_trigger_edge_state,trigger_edge_state}==2'b10)
            trigger_edge_o<=!trigger_edge_o;
        else
            trigger_edge_o<=trigger_edge_o;
    end
    //���л������λ�������
    wire h_exceed;
    wire v_exceed;
    assign h_exceed = I_vtc2_offset_x + H2_ActiveSize > H_Visible_area - 1'b1;
    assign v_exceed = I_vtc2_offset_y + V2_ActiveSize > V_Visible_area - 1'b1;
    assign hs2_valid = h_exceed ? (visible_hcount >= I_vtc2_offset_x && visible_hcount < H_Visible_area):
                                  (visible_hcount >= I_vtc2_offset_x && visible_hcount < I_vtc2_offset_x + H2_ActiveSize);  
  
    assign vs2_valid = v_exceed ? (visible_vcount >= I_vtc2_offset_y && visible_vcount < V_Visible_area):
                                  (visible_vcount >= I_vtc2_offset_y && visible_vcount < I_vtc2_offset_y + V2_ActiveSize);
  
    wire vtc2_de    =  hs2_valid && vs2_valid; //���л���������Ч�����ź�
    reg   O_vtc2_de;
    reg [2:0]rst_cnt;
    /*reg [4:0]frame_cnt;
    always @(posedge clk_ctrl or negedge reset_n)begin //ͨ������������ͬ����λ
       if(reset_n == 1'b0)
           frame_cnt <= 5'b11111;
        else if(Frame_Begin)
            frame_cnt<=5'b00000;
       else if(frame_cnt[4] == 1'b0)
           frame_cnt <= frame_cnt + 1'b1;
   end    
    wire frame_rst=(frame_cnt==5'b00000)?0:1;*/
    always @(posedge clk_ctrl or negedge reset_n)begin //ͨ������������ͬ����λ
       if(reset_n == 1'b0)
           rst_cnt <= 3'd0;
       else if(rst_cnt[2] == 1'b0)
           rst_cnt <= rst_cnt + 1'b1;
   end    
    wire rst_sync = rst_cnt[2]; //ͬ����λ   
    //��һ�μĴ��������������ڸ���ʱ��������ڸ߷ֱ��ʣ����ٵ��źţ����Ŀ��Ը����ڲ�ʱ���������ڸ����ٶ�
    always @(posedge clk_ctrl)begin
        if(rst_sync == 1'b0)begin
            O_vtc_vs <= 1'b0;
            O_vtc_hs <= 1'b0;
            O_vtc_de <= 1'b0;
            O_vtc2_de <= 1'b0;
        end
        else begin
            O_vtc_vs <= I_vtc_vs; //��ͬ���źŴ������
            O_vtc_hs <= I_vtc_hs; //��ͬ���źŴ������
            O_vtc_de <= I_vtc_de; //��Ƶ��Ч�źŴ������
            O_vtc2_de <= vtc2_de; //���л���������Ч�����ź�
        end
    end
    
    uiwave uiwave
    (
    //����1
    .I_wave1_clk(I_wave1_clk),      //����1ʱ��
    .I_wave1_data(I_wave1_data),     //����1����
    .I_wave1_data_de(I_wave1_data_de),  //����1������Ч
    
    //����2
    .I_wave2_clk(I_wave2_clk),      //����2ʱ��
    .I_wave2_data(I_wave2_data),     //����2����
    .I_wave2_data_de(I_wave2_data_de),  //����2������Ч
    
    //VTCʱ������
    .I_vtc_rstn(reset_n),       //ʱ��λ����
    .I_vtc_clk(clk_ctrl),        //ʱ��ʱ������
    .I_vtc_vs(O_vtc_vs),         //VS-֡ͬ�����ź�ͬ������
    .I_vtc_de(O_vtc2_de),         //de��Ч�����ź�ͬ������
    
    //ͬ��ʱ��������Լ��������
    .O_vtc_vs(),         //֡ͬ�����
    .O_vtc_de(),         //de�ź�ͬ�������
    .O_vtc_rgb(O_vtc_rgb),     //ͬ�������ʾ��ɫ

    .single_flag(single_flag),
    .trigger_edge(trigger_edge_o),
    .trigger_button_flag(trigger_button_minus_flag)
    );
endmodule