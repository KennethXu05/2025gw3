//Copyright (C)2014-2025 Gowin Semiconductor Corporation.
//All rights reserved.
//File Title: IP file
//Tool Version: V1.9.12 (64-bit)
//Part Number: GW5AT-LV138PG484AC1/I0
//Device: GW5AT-138
//Device Version: B
//Created Time: Mon Oct 13 16:24:36 2025

module asscii_rom (dout, clk, oce, ce, reset, ad);

output [15:0] dout;
input clk;
input oce;
input ce;
input reset;
input [11:0] ad;

wire lut_f_0;
wire lut_f_1;
wire [23:0] prom_inst_0_dout_w;
wire [7:0] prom_inst_0_dout;
wire [23:0] prom_inst_1_dout_w;
wire [15:8] prom_inst_1_dout;
wire [15:0] prom_inst_2_dout_w;
wire [15:0] prom_inst_2_dout;
wire dff_q_0;
wire gw_gnd;

assign gw_gnd = 1'b0;

LUT2 lut_inst_0 (
  .F(lut_f_0),
  .I0(ce),
  .I1(ad[11])
);
defparam lut_inst_0.INIT = 4'h2;
LUT3 lut_inst_1 (
  .F(lut_f_1),
  .I0(ce),
  .I1(ad[10]),
  .I2(ad[11])
);
defparam lut_inst_1.INIT = 8'h20;
pROM prom_inst_0 (
    .DO({prom_inst_0_dout_w[23:0],prom_inst_0_dout[7:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_0),
    .RESET(reset),
    .AD({ad[10:0],gw_gnd,gw_gnd,gw_gnd})
);

defparam prom_inst_0.READ_MODE = 1'b0;
defparam prom_inst_0.BIT_WIDTH = 8;
defparam prom_inst_0.RESET_MODE = "SYNC";
defparam prom_inst_0.INIT_RAM_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_01 = 256'h0000000080C0C0800000008080808080808080C0C0C0C0C0C0C0000000000000;
defparam prom_inst_0.INIT_RAM_02 = 256'h000000000000000000000000000000000000000000000080C060703838180000;
defparam prom_inst_0.INIT_RAM_03 = 256'h000000002020202030FEFEFE101010101010FEFEFE0808080808000000000000;
defparam prom_inst_0.INIT_RAM_04 = 256'h00000000C06030181818183830F0E0C0000000003838181830C0000000000000;
defparam prom_inst_0.INIT_RAM_05 = 256'h00000000386C44C6C6C6C6C6C6446C3880808040404020201010000000000000;
defparam prom_inst_0.INIT_RAM_06 = 256'h00000000387CE6C2C02020201010107C00000000808080800000000000000000;
defparam prom_inst_0.INIT_RAM_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_08 = 256'h000204081830206040C0C0808080808080808080C0C040602030180804020000;
defparam prom_inst_0.INIT_RAM_09 = 256'h0000000000000000000000808080808080808080000000000000000000000000;
defparam prom_inst_0.INIT_RAM_0A = 256'h0000000000000000C0C0C0868E9CB0C0C0B09C8EC6C0C0C00000000000000000;
defparam prom_inst_0.INIT_RAM_0B = 256'h000000000000000080808080808080FE80808080808080000000000000000000;
defparam prom_inst_0.INIT_RAM_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_0D = 256'h000000000000000000000000000000FE00000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_0F = 256'h0000000000000000000000000000008080C0406020301018080C040602000000;
defparam prom_inst_0.INIT_RAM_10 = 256'h00000000C020301818080C0C0C0C0C0C0C0C0C0C0818183020C0000000000000;
defparam prom_inst_0.INIT_RAM_11 = 256'h00000000F8C08080808080808080808080808080808080808080000000000000;
defparam prom_inst_0.INIT_RAM_12 = 256'h00000000F8F80C040404000080C0603018180C0C0C0C0C1838E0000000000000;
defparam prom_inst_0.INIT_RAM_13 = 256'h00000000C03018080C0C0C0C081870C0603018181818183060C0000000000000;
defparam prom_inst_0.INIT_RAM_14 = 256'h00000000FC6060606060FC6060606060606060606060E0E06060000000000000;
defparam prom_inst_0.INIT_RAM_15 = 256'h00000000C03018180C0C0C0C0C0C081830E0000000000000FCFC000000000000;
defparam prom_inst_0.INIT_RAM_16 = 256'h00000000E03018080C0C0C0C0C0C081830E000000000181818E0000000000000;
defparam prom_inst_0.INIT_RAM_17 = 256'h000000000000000000000000000080804040402020101008FCFC000000000000;
defparam prom_inst_0.INIT_RAM_18 = 256'h00000000C030180C0C0C0C1C3878F0C02018080C0C0C0C1830E0000000000000;
defparam prom_inst_0.INIT_RAM_19 = 256'h0000000080C060301018180C8C6C2C1C0C0C0C0C0C08181020C0000000000000;
defparam prom_inst_0.INIT_RAM_1A = 256'h0000000080C0C0800000000000000080C0C08000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_1B = 256'h0000008080808000000000000000008080800000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_1C = 256'h0000000004081020408000000000000000000000804020100804000000000000;
defparam prom_inst_0.INIT_RAM_1D = 256'h000000000000000000000000FE0000000000FE00000000000000000000000000;
defparam prom_inst_0.INIT_RAM_1E = 256'h0000000000000000000080402010080810204080000000000000000000000000;
defparam prom_inst_0.INIT_RAM_1F = 256'h0000000080C0C080000080808080C070180C06060606060C18E0000000000000;
defparam prom_inst_0.INIT_RAM_20 = 256'h00000000E0180C040230E8646462222222223232B2D4040810E0000000000000;
defparam prom_inst_0.INIT_RAM_21 = 256'h000000003E1C181818303030F02060606040C0C0C0C080808080000000000000;
defparam prom_inst_0.INIT_RAM_22 = 256'h00000000F0180C0606060606040C18E030180C0C0C0C0C1838E0000000000000;
defparam prom_inst_0.INIT_RAM_23 = 256'h00000000E01008040202000000000000000000000202060C1CE0000000000000;
defparam prom_inst_0.INIT_RAM_24 = 256'h00000000C06018180C0C040606060606060606060C0C081870C0000000000000;
defparam prom_inst_0.INIT_RAM_25 = 256'h00000000FC0C040202000000101030F030101000000202040CFC000000000000;
defparam prom_inst_0.INIT_RAM_26 = 256'h000000000000000000000010101030F030101000000202041CFC000000000000;
defparam prom_inst_0.INIT_RAM_27 = 256'h00000000C020181818181818187E0000000000000808181030C0000000000000;
defparam prom_inst_0.INIT_RAM_28 = 256'h000000003F0C0C0C0C0C0C0C0C0C0CFC0C0C0C0C0C0C0C0C0C3F000000000000;
defparam prom_inst_0.INIT_RAM_29 = 256'h00000000F88080808080808080808080808080808080808080F8000000000000;
defparam prom_inst_0.INIT_RAM_2A = 256'h0080C060606060606060606060606060606060606060606060FE000000000000;
defparam prom_inst_0.INIT_RAM_2B = 256'h000000003E18183030306060C0C080800000008080406020307C000000000000;
defparam prom_inst_0.INIT_RAM_2C = 256'h00000000FC0C0402020000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_2D = 256'h000000003F0C0C0C8C8C8C8C4C4C4C4C4C2C2C2C2C1C1C1C1C0F000000000000;
defparam prom_inst_0.INIT_RAM_2E = 256'h00000000040C0C1C1C34346464C4C4848404040404040404041F000000000000;
defparam prom_inst_0.INIT_RAM_2F = 256'h00000000C03018080C0C060606060606060606040C0C081830C0000000000000;
defparam prom_inst_0.INIT_RAM_30 = 256'h0000000000000000000000000000E0180C0606060606060C18F0000000000000;
defparam prom_inst_0.INIT_RAM_31 = 256'h001C3C32E070786CCC84060606060606060606060C0C081830C0000000000000;
defparam prom_inst_0.INIT_RAM_32 = 256'h000000001E1818303030606060C0C0E030180C0C0C0C0C1838E0000000000000;
defparam prom_inst_0.INIT_RAM_33 = 256'h00000000E030180C0C0C0C1C1878F0C0000000000808181878C8000000000000;
defparam prom_inst_0.INIT_RAM_34 = 256'h00000000E08080808080808080808080808080808082828684FC000000000000;
defparam prom_inst_0.INIT_RAM_35 = 256'h00000000C020100808080808080808080808080808080808083E000000000000;
defparam prom_inst_0.INIT_RAM_36 = 256'h0000000000008080804040404020202020101010100808080C1E000000000000;
defparam prom_inst_0.INIT_RAM_37 = 256'h000000002020203070707070686848C8C8C8C4C4C484848486CF000000000000;
defparam prom_inst_0.INIT_RAM_38 = 256'h000000003E1C183030706060C0C080808080404020201010083E000000000000;
defparam prom_inst_0.INIT_RAM_39 = 256'h00000000E080808080808080808080404020202010101008083E000000000000;
defparam prom_inst_0.INIT_RAM_3A = 256'h00000000FC1C04060200000000008080C0C060603018180C0CFE000000000000;
defparam prom_inst_0.INIT_RAM_3B = 256'h0000FC00000000000000000000000000000000000000000000000000FC000000;
defparam prom_inst_0.INIT_RAM_3C = 256'h00060C0C0C1818303030606040C0808080000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_3D = 256'h0000C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0C0000000;
defparam prom_inst_0.INIT_RAM_3E = 256'h00000000000000000000000000000000000000000000000000001020E0C00000;
defparam prom_inst_0.INIT_RAM_3F = 256'hFF00000000000000000000000000000000000000000000000000000000000000;

pROM prom_inst_1 (
    .DO({prom_inst_1_dout_w[23:0],prom_inst_1_dout[15:8]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_0),
    .RESET(reset),
    .AD({ad[10:0],gw_gnd,gw_gnd,gw_gnd})
);

defparam prom_inst_1.READ_MODE = 1'b0;
defparam prom_inst_1.BIT_WIDTH = 8;
defparam prom_inst_1.RESET_MODE = "SYNC";
defparam prom_inst_1.INIT_RAM_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_1.INIT_RAM_01 = 256'h0000000001030301000000010101010101010101030303030303000000000000;
defparam prom_inst_1.INIT_RAM_02 = 256'h000000000000000000000000000000000000000000002131180C0E0707030000;
defparam prom_inst_1.INIT_RAM_03 = 256'h0000000010101010187F7F7F0808080808087F7F7F0404040404000000000000;
defparam prom_inst_1.INIT_RAM_04 = 256'h00010101071931313939010101010103070F0D1D191919090D03010100000000;
defparam prom_inst_1.INIT_RAM_05 = 256'h0000000010100808080404020202396D44C6C6C6C6C6C6446C38000000000000;
defparam prom_inst_1.INIT_RAM_06 = 256'h000000001E3160C1C1C3C7C6CE4C3C381C3A333131313131190F000000000000;
defparam prom_inst_1.INIT_RAM_07 = 256'h000000000000000000000000000000000000000000006030080C0C3C3C380000;
defparam prom_inst_1.INIT_RAM_08 = 256'h0000000000000000000000010101010101010101000000000000000000000000;
defparam prom_inst_1.INIT_RAM_09 = 256'h00402010180C040603030301010101010101010103030206040C181020400000;
defparam prom_inst_1.INIT_RAM_0A = 256'h000000000000000001010131381C060101061C38300101000000000000000000;
defparam prom_inst_1.INIT_RAM_0B = 256'h0000000000000000000000000000003F00000000000000000000000000000000;
defparam prom_inst_1.INIT_RAM_0C = 256'h6030080C0C3C3C38000000000000000000000000000000000000000000000000;
defparam prom_inst_1.INIT_RAM_0D = 256'h0000000000000000000000000000007F00000000000000000000000000000000;
defparam prom_inst_1.INIT_RAM_0E = 256'h00000000183C3C18000000000000000000000000000000000000000000000000;
defparam prom_inst_1.INIT_RAM_0F = 256'h0000406020301018080C04060203010100000000000000000000000000000000;
defparam prom_inst_1.INIT_RAM_10 = 256'h0000000003060C181818303030303030303030301818180C0603000000000000;
defparam prom_inst_1.INIT_RAM_11 = 256'h000000001F0301010101010101010101010101010101011F0100000000000000;
defparam prom_inst_1.INIT_RAM_12 = 256'h000000003F3F2010080402030100000000000030302020100807000000000000;
defparam prom_inst_1.INIT_RAM_13 = 256'h0000000007183030303000000000000300000000303030301807000000000000;
defparam prom_inst_1.INIT_RAM_14 = 256'h000000000300000000007F402030100808040402010100000000000000000000;
defparam prom_inst_1.INIT_RAM_15 = 256'h0000000007182020303000000000101814131010101010100F0F000000000000;
defparam prom_inst_1.INIT_RAM_16 = 256'h00000000030E0C181830303030303838363330101018080C0601000000000000;
defparam prom_inst_1.INIT_RAM_17 = 256'h0000000003030303030301010101000000000000202030101F1F000000000000;
defparam prom_inst_1.INIT_RAM_18 = 256'h000000000718306060606060303018070F1E3838303030180C07000000000000;
defparam prom_inst_1.INIT_RAM_19 = 256'h000000000F303030000000000F18307060606060606030301807000000000000;
defparam prom_inst_1.INIT_RAM_1A = 256'h0000000001030301000000000000000103030100000000000000000000000000;
defparam prom_inst_1.INIT_RAM_1B = 256'h0003030103030300000000000000000303030000000000000000000000000000;
defparam prom_inst_1.INIT_RAM_1C = 256'h0000000000000000000001020408101008040201000000000000000000000000;
defparam prom_inst_1.INIT_RAM_1D = 256'h0000000000000000000000007F00000000007F00000000000000000000000000;
defparam prom_inst_1.INIT_RAM_1E = 256'h0000000020100804020100000000000000000000010204081020000000000000;
defparam prom_inst_1.INIT_RAM_1F = 256'h0000000001030301000000000000000000003838383010180C03000000000000;
defparam prom_inst_1.INIT_RAM_20 = 256'h00000000030C18103033266666666666666363213130180C0603000000000000;
defparam prom_inst_1.INIT_RAM_21 = 256'h00000000F8602020201010101F180808080C0404040403030303000000000000;
defparam prom_inst_1.INIT_RAM_22 = 256'h000000007F181818181818181818181F1818181818181818187F000000000000;
defparam prom_inst_1.INIT_RAM_23 = 256'h00000000030C1810303060606060606060606030303018080603000000000000;
defparam prom_inst_1.INIT_RAM_24 = 256'h000000007F18181818181818181818181818181818181818187F000000000000;
defparam prom_inst_1.INIT_RAM_25 = 256'h000000007F181818181818181818181F1818181818181818187F000000000000;
defparam prom_inst_1.INIT_RAM_26 = 256'h000000007E181818181818181818181F1818181818181818187F000000000000;
defparam prom_inst_1.INIT_RAM_27 = 256'h00000000070C1810303020606060606060606020303018080C03000000000000;
defparam prom_inst_1.INIT_RAM_28 = 256'h00000000FC303030303030303030303F303030303030303030FC000000000000;
defparam prom_inst_1.INIT_RAM_29 = 256'h000000001F01010101010101010101010101010101010101011F000000000000;
defparam prom_inst_1.INIT_RAM_2A = 256'h3F71707000000000000000000000000000000000000000000007000000000000;
defparam prom_inst_1.INIT_RAM_2B = 256'h000000007E1818181818181818181D1D1B19191818181818187E000000000000;
defparam prom_inst_1.INIT_RAM_2C = 256'h000000007F18181818181818181818181818181818181818187E000000000000;
defparam prom_inst_1.INIT_RAM_2D = 256'h00000000F1212323232322262626262C2C2C2C2C3838383838F0000000000000;
defparam prom_inst_1.INIT_RAM_2E = 256'h00000000F8202020202020202020202121232326262C2C3838F0000000000000;
defparam prom_inst_1.INIT_RAM_2F = 256'h00000000030C1810303020606060606060606060303010180C03000000000000;
defparam prom_inst_1.INIT_RAM_30 = 256'h000000007E1818181818181818181F181818181818181818187F000000000000;
defparam prom_inst_1.INIT_RAM_31 = 256'h00000000030C1838382760606060606060606060303010180C03000000000000;
defparam prom_inst_1.INIT_RAM_32 = 256'h000000007E181818181818181818181F1818181818181818187F000000000000;
defparam prom_inst_1.INIT_RAM_33 = 256'h000000002738302060404000000001071F3C706060606030180F000000000000;
defparam prom_inst_1.INIT_RAM_34 = 256'h000000000701010101010101010101010101010101414121313F000000000000;
defparam prom_inst_1.INIT_RAM_35 = 256'h00000000071C18303030303030303030303030303030303030FC000000000000;
defparam prom_inst_1.INIT_RAM_36 = 256'h000000000101010103030303060606060C0C0C0C0C181818187C000000000000;
defparam prom_inst_1.INIT_RAM_37 = 256'h0000000008080C0C0C0C1C1A1A1A1211313131313020216161F3000000000000;
defparam prom_inst_1.INIT_RAM_38 = 256'h000000007C101808080404020201010101030306060C0C18187C000000000000;
defparam prom_inst_1.INIT_RAM_39 = 256'h000000000701010101010101010103030306060C0C0C1818387E000000000000;
defparam prom_inst_1.INIT_RAM_3A = 256'h000000007F303018180C06060303010100000000002030181C1F000000000000;
defparam prom_inst_1.INIT_RAM_3B = 256'h0000030303030303030303030303030303030303030303030303030303000000;
defparam prom_inst_1.INIT_RAM_3C = 256'h00000000000000000000000000000001010103020606040C0818180000000000;
defparam prom_inst_1.INIT_RAM_3D = 256'h00003F000000000000000000000000000000000000000000000000003F000000;
defparam prom_inst_1.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000080603030000;
defparam prom_inst_1.INIT_RAM_3F = 256'hFF00000000000000000000000000000000000000000000000000000000000000;

pROM prom_inst_2 (
    .DO({prom_inst_2_dout_w[15:0],prom_inst_2_dout[15:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_1),
    .RESET(reset),
    .AD({ad[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam prom_inst_2.READ_MODE = 1'b0;
defparam prom_inst_2.BIT_WIDTH = 16;
defparam prom_inst_2.RESET_MODE = "SYNC";
defparam prom_inst_2.INIT_RAM_00 = 256'h00000000000000000000000000000000000000000000008003001E0000000000;
defparam prom_inst_2.INIT_RAM_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_2.INIT_RAM_02 = 256'h3018183007E00000000000000000000000000000000000000000000000000000;
defparam prom_inst_2.INIT_RAM_03 = 256'h00000000000000001F8E3079601960186018601830181C1807D8003830183018;
defparam prom_inst_2.INIT_RAM_04 = 256'h1C181A3819E01800180018001800180018007800080000000000000000000000;
defparam prom_inst_2.INIT_RAM_05 = 256'h000000000000000013E01C301C181808180C180C180C180C180C180C180C1C0C;
defparam prom_inst_2.INIT_RAM_06 = 256'h0C180E1003E00000000000000000000000000000000000000000000000000000;
defparam prom_inst_2.INIT_RAM_07 = 256'h000000000000000003E00C101808180430043000300030003000300030181818;
defparam prom_inst_2.INIT_RAM_08 = 256'h18180C3807D80018001800180018001800180078000800000000000000000000;
defparam prom_inst_2.INIT_RAM_09 = 256'h000000000000000007900C5E1838101830183018301830183018301830181818;
defparam prom_inst_2.INIT_RAM_0A = 256'h08180C3003C00000000000000000000000000000000000000000000000000000;
defparam prom_inst_2.INIT_RAM_0B = 256'h000000000000000003E00E18180818043000300030003FFC300C300C300C1808;
defparam prom_inst_2.INIT_RAM_0C = 256'h030003003FF8030003000300030601060186007C000000000000000000000000;
defparam prom_inst_2.INIT_RAM_0D = 256'h00000000000000001FF003000300030003000300030003000300030003000300;
defparam prom_inst_2.INIT_RAM_0E = 256'h08180C3603EE0000000000000000000000000000000000000000000000000000;
defparam prom_inst_2.INIT_RAM_0F = 256'h07E01818300C300C300C181C0FF81FC0180018000FE00C300818181818181818;
defparam prom_inst_2.INIT_RAM_10 = 256'h1C181A3019E01800180018001800180018007800080000000000000000000000;
defparam prom_inst_2.INIT_RAM_11 = 256'h00000000000000007E7E18181818181818181818181818181818181818181818;
defparam prom_inst_2.INIT_RAM_12 = 256'h018001801F800080000000000000018003C00180000000000000000000000000;
defparam prom_inst_2.INIT_RAM_13 = 256'h00000000000000001FF801800180018001800180018001800180018001800180;
defparam prom_inst_2.INIT_RAM_14 = 256'h0030003003F00010000000000000003000780038000000000000000000000000;
defparam prom_inst_2.INIT_RAM_15 = 256'h0F80184018600030003000300030003000300030003000300030003000300030;
defparam prom_inst_2.INIT_RAM_16 = 256'h18201830187C1800180018001800180018007800080000000000000000000000;
defparam prom_inst_2.INIT_RAM_17 = 256'h00000000000000007E3E181C18181830183018601CC01EC01B80198018801840;
defparam prom_inst_2.INIT_RAM_18 = 256'h0180018001800180018001800180018001801F80008000000000000000000000;
defparam prom_inst_2.INIT_RAM_19 = 256'h00000000000000001FF801800180018001800180018001800180018001800180;
defparam prom_inst_2.INIT_RAM_1A = 256'h618671C6EF3C2000000000000000000000000000000000000000000000000000;
defparam prom_inst_2.INIT_RAM_1B = 256'h0000000000000000F3CF61866186618661866186618661866186618661866186;
defparam prom_inst_2.INIT_RAM_1C = 256'h1C187A3009E00000000000000000000000000000000000000000000000000000;
defparam prom_inst_2.INIT_RAM_1D = 256'h00000000000000007E7E18181818181818181818181818181818181818181818;
defparam prom_inst_2.INIT_RAM_1E = 256'h08180C3003C00000000000000000000000000000000000000000000000000000;
defparam prom_inst_2.INIT_RAM_1F = 256'h000000000000000003C00C3018181818300C300C300C300C300C300C100C1818;
defparam prom_inst_2.INIT_RAM_20 = 256'h1C187A3009E00000000000000000000000000000000000000000000000000000;
defparam prom_inst_2.INIT_RAM_21 = 256'h7E0018001800180019E01E301C181818180C180C180C180C180C180C180C1808;
defparam prom_inst_2.INIT_RAM_22 = 256'h18380C7803C80000000000000000000000000000000000000000000000000000;
defparam prom_inst_2.INIT_RAM_23 = 256'h007E00180018001807980C781838101830183018301830183018301830181818;
defparam prom_inst_2.INIT_RAM_24 = 256'h06867E66061C0000000000000000000000000000000000000000000000000000;
defparam prom_inst_2.INIT_RAM_25 = 256'h00000000000000007FE006000600060006000600060006000600060007000780;
defparam prom_inst_2.INIT_RAM_26 = 256'h0C0C061C03E40000000000000000000000000000000000000000000000000000;
defparam prom_inst_2.INIT_RAM_27 = 256'h000000000000000013F01C18180C100C100C001C007801F007C00E000C040C04;
defparam prom_inst_2.INIT_RAM_28 = 256'h030003003FF80700030001000100010000000000000000000000000000000000;
defparam prom_inst_2.INIT_RAM_29 = 256'h000000000000000000F001880304030403000300030003000300030003000300;
defparam prom_inst_2.INIT_RAM_2A = 256'h1818181878780808000000000000000000000000000000000000000000000000;
defparam prom_inst_2.INIT_RAM_2B = 256'h000000000000000007900C5E1838181818181818181818181818181818181818;
defparam prom_inst_2.INIT_RAM_2C = 256'h1808180C7C3E0000000000000000000000000000000000000000000000000000;
defparam prom_inst_2.INIT_RAM_2D = 256'h000000000000000001000180018003C0034003400620062004200C100C101818;
defparam prom_inst_2.INIT_RAM_2E = 256'h21846186FBCF0000000000000000000000000000000000000000000000000000;
defparam prom_inst_2.INIT_RAM_2F = 256'h000000000000000004200C200C300C700E701A701A481AC811C831C831843184;
defparam prom_inst_2.INIT_RAM_30 = 256'h0E100C103E7C0000000000000000000000000000000000000000000000000000;
defparam prom_inst_2.INIT_RAM_31 = 256'h00000000000000007C7E1818081804300460026001C001800180034003400620;
defparam prom_inst_2.INIT_RAM_32 = 256'h181018187C3E0000000000000000000000000000000000000000000000000000;
defparam prom_inst_2.INIT_RAM_33 = 256'h3C003E000200010001000100018001800140034002400620062004200C100810;
defparam prom_inst_2.INIT_RAM_34 = 256'h303030383FF80000000000000000000000000000000000000000000000000000;
defparam prom_inst_2.INIT_RAM_35 = 256'h00000000000000003FF83018180C0C040E04060003000380018000C020E02060;
defparam prom_inst_2.INIT_RAM_36 = 256'h00C0002000200020002000200020002000200020002000200010000C00000000;
defparam prom_inst_2.INIT_RAM_37 = 256'h0000000C00100020002000200020002000200020002000200020002000400180;
defparam prom_inst_2.INIT_RAM_38 = 256'h0080008000800080008000800080008000800080008000800080008000800080;
defparam prom_inst_2.INIT_RAM_39 = 256'h0080008000800080008000800080008000800080008000800080008000800080;
defparam prom_inst_2.INIT_RAM_3A = 256'h0180020002000200020002000200020002000200020002000400180000000000;
defparam prom_inst_2.INIT_RAM_3B = 256'h00001800040002000200020002000200020002000200020002000200010000C0;
defparam prom_inst_2.INIT_RAM_3C = 256'h000000000000000000000000000000000000003800E44082418223001E000000;
defparam prom_inst_2.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;

DFFRE dff_inst_0 (
  .Q(dff_q_0),
  .D(ad[11]),
  .CLK(clk),
  .CE(ce),
  .RESET(gw_gnd)
);
MUX2 mux_inst_2 (
  .O(dout[0]),
  .I0(prom_inst_0_dout[0]),
  .I1(prom_inst_2_dout[0]),
  .S0(dff_q_0)
);
MUX2 mux_inst_5 (
  .O(dout[1]),
  .I0(prom_inst_0_dout[1]),
  .I1(prom_inst_2_dout[1]),
  .S0(dff_q_0)
);
MUX2 mux_inst_8 (
  .O(dout[2]),
  .I0(prom_inst_0_dout[2]),
  .I1(prom_inst_2_dout[2]),
  .S0(dff_q_0)
);
MUX2 mux_inst_11 (
  .O(dout[3]),
  .I0(prom_inst_0_dout[3]),
  .I1(prom_inst_2_dout[3]),
  .S0(dff_q_0)
);
MUX2 mux_inst_14 (
  .O(dout[4]),
  .I0(prom_inst_0_dout[4]),
  .I1(prom_inst_2_dout[4]),
  .S0(dff_q_0)
);
MUX2 mux_inst_17 (
  .O(dout[5]),
  .I0(prom_inst_0_dout[5]),
  .I1(prom_inst_2_dout[5]),
  .S0(dff_q_0)
);
MUX2 mux_inst_20 (
  .O(dout[6]),
  .I0(prom_inst_0_dout[6]),
  .I1(prom_inst_2_dout[6]),
  .S0(dff_q_0)
);
MUX2 mux_inst_23 (
  .O(dout[7]),
  .I0(prom_inst_0_dout[7]),
  .I1(prom_inst_2_dout[7]),
  .S0(dff_q_0)
);
MUX2 mux_inst_26 (
  .O(dout[8]),
  .I0(prom_inst_1_dout[8]),
  .I1(prom_inst_2_dout[8]),
  .S0(dff_q_0)
);
MUX2 mux_inst_29 (
  .O(dout[9]),
  .I0(prom_inst_1_dout[9]),
  .I1(prom_inst_2_dout[9]),
  .S0(dff_q_0)
);
MUX2 mux_inst_32 (
  .O(dout[10]),
  .I0(prom_inst_1_dout[10]),
  .I1(prom_inst_2_dout[10]),
  .S0(dff_q_0)
);
MUX2 mux_inst_35 (
  .O(dout[11]),
  .I0(prom_inst_1_dout[11]),
  .I1(prom_inst_2_dout[11]),
  .S0(dff_q_0)
);
MUX2 mux_inst_38 (
  .O(dout[12]),
  .I0(prom_inst_1_dout[12]),
  .I1(prom_inst_2_dout[12]),
  .S0(dff_q_0)
);
MUX2 mux_inst_41 (
  .O(dout[13]),
  .I0(prom_inst_1_dout[13]),
  .I1(prom_inst_2_dout[13]),
  .S0(dff_q_0)
);
MUX2 mux_inst_44 (
  .O(dout[14]),
  .I0(prom_inst_1_dout[14]),
  .I1(prom_inst_2_dout[14]),
  .S0(dff_q_0)
);
MUX2 mux_inst_47 (
  .O(dout[15]),
  .I0(prom_inst_1_dout[15]),
  .I1(prom_inst_2_dout[15]),
  .S0(dff_q_0)
);
endmodule //asscii_rom
