
 module uiwave
 (
 //����1
 input         I_wave1_clk,      //����1ʱ��
 input  [7 :0] I_wave1_data,     //����1����
 input         I_wave1_data_de,  //����1������Ч
 
 //����2
 input         I_wave2_clk,      //����2ʱ��
 input  [7 :0] I_wave2_data,     //����2����
 input         I_wave2_data_de,  //����2������Ч
 
 //VTCʱ������
 input         I_vtc_rstn,       //ʱ��λ����
 input         I_vtc_clk,        //ʱ��ʱ������
 input         I_vtc_vs,         //VS-֡ͬ�����ź�ͬ������
 input         I_vtc_de,         //de��Ч�����ź�ͬ������
 
 //ͬ��ʱ��������Լ��������
 output        O_vtc_vs,         //֡ͬ�����
 output        O_vtc_de,         //de�ź�ͬ�������
 output reg [15:0] O_vtc_rgb,     //ͬ�������ʾ��ɫ
 input         single_flag,


 input trigger_edge,
 input trigger_button_flag
 );
 
 reg  [1 :0] vtc_vs_r; //vs�Ĵ���
 reg  [1 :0] vtc_de_r; //de�Ĵ���
 reg  [11 :0] vcnt,hcnt;//vcnt�����ж����У�hcnt�����ж�����
 
 reg    grid_de; //դ�����ʹ��
 
 assign O_vtc_vs = vtc_vs_r[0]; //ͬ�������O_vtc_vs
 assign O_vtc_de = vtc_de_r[0]; //ͬ�������O_vtc_de
 
 //�Ĵ�,ͬ��
 always @(posedge I_vtc_clk)begin
     vtc_vs_r <= {vtc_vs_r[0],I_vtc_vs};
     vtc_de_r <= {vtc_de_r[0],I_vtc_de};
 end
 /*
 reg [27:0]trigger_cnt;
 always @(posedge I_vtc_clk or negedge I_vtc_rstn) begin
    if(I_vtc_rstn==0)
        trigger_cnt<=0;
    else if(trigger_button_flag)
        trigger_cnt<=trigger_cnt+1;
    else if(trigger_cnt>=28'd199_999_999)
        trigger_cnt<=0;
    else
        trigger_cnt<=0;
 end*/
 //����hcnt���ڼ����У�vcnt���ڼ�������
 
 //hcnt���ؼ�����
 always @(posedge I_vtc_clk)begin
     if(hcnt == 749)
         hcnt <= 12'd0;
     else if(vtc_de_r[0] && (hcnt != 749)) //hcnt�����У�����512������
         hcnt <= hcnt + 1'b1;
 end
 
 //vcnt�����ж�����
 always @(posedge I_vtc_clk)begin
     if(vtc_vs_r == 2'b01)
         vcnt <= 12'd0;
     else if((vtc_de_r == 2'b10) && (vcnt != 255)) //��de�ź����ڼ����У�����256��
         vcnt <= vcnt + 1'b1;
 end
 
 //դ�����
   /*  wire h_grid = (hcnt[2:0] == 3'd7) && (vcnt[5:0] == 6'd63 || vcnt == 10'd0);
    // ����2������դ���ߣ����ߣ�
    // ÿ64�У�0��64��128...608�������ڵ�7�У�ÿ8��1���㣩
    wire v_grid = (vcnt[2:0] == 3'd7) && (hcnt[5:0] == 6'd63 || hcnt == 10'd0);
    // ����3��ԭ���ǣ�0,0��
    wire origin = (hcnt == 10'd0) && (vcnt == 10'd0);
    
 // դ����ƣ�����640��480��Ч��ʾ����

always @(posedge I_vtc_clk) begin
    // ����1������դ���ߣ����ߣ�
    // ÿ64�У�0��64��128...448�������ڵ�7�У�ÿ8��1���㣩

    // դ����Ч�źţ�������һ������������ʾ��Ч������
    grid_de <= (h_grid || v_grid || origin) && O_vtc_de;
end*/
reg [7:0]trigger_line;
reg trigger_de;
always @(posedge I_vtc_clk or negedge I_vtc_rstn) begin
    if(I_vtc_rstn==1'b0)
        trigger_line<=8'h00;
    else if(trigger_button_flag)
        trigger_line<=trigger_line+1'b1;
    else
        trigger_line<=trigger_line;
end

 always @(posedge I_vtc_clk)begin
     if((hcnt[2:0]==7&&(vcnt[5:0]==63||vcnt == 0))||((hcnt[5:0]==63||hcnt==0)&&vcnt[2:0]==7)||(vcnt == 0 && hcnt==0)) 
         grid_de <= O_vtc_de;
     else 
         grid_de <= 1'b0;
 end 
 always @(posedge I_vtc_clk)begin
     if(hcnt[1:0]==3&&vcnt[7:0]==trigger_line) 
         trigger_de <= O_vtc_de;
     else 
         trigger_de <= 1'b0;
 end 
 //1--���Ʋ�������1����ɫ��
 //2--���Ʋ�������2����ɫ��
 //3--����դ�����ߣ���ɫ��
 //4--���Ʊ���ɫ����ɫ
 always @(posedge I_vtc_clk)begin
     casex({grid_de,trigger_de,wave1_pixel_en})
             3'bxx1:
                O_vtc_rgb <= {5'b00000,6'b111111,5'b00000};   //wave1�ź���ʾ������ɫ
             3'bx10:
                O_vtc_rgb <= {5'b11111,6'b000000,5'b11111};   //������ʾ����Ϊ��ɫ��
             3'b100:
                O_vtc_rgb <= {5'b10010,6'b100101,5'b10010};   //������ʾ����Ϊ��ɫ��
         default:
                O_vtc_rgb <= {5'b00000,6'b000000,5'b00000};   //��ɫ����
     endcase
 end 
 
 //���λ���1���Լ����λ������ص����ʹ��
 uiwave_buf uiwave1_buf_inst
 (
 .I_wave_clk(I_wave1_clk),  //д��������ʱ�ӣ���ADC�ɼ�ʱ��ͬ��
 .I_wave_data(I_wave1_data),//д����
 .I_wave_data_de(I_wave1_data_de),//д������Ч
 .I_vtc_clk(I_vtc_clk),    //VTCʱ������ʱ������
 .I_vtc_rstn(I_vtc_rstn),  //VTCʱ��������λ 
 .I_vtc_de_r(vtc_de_r[0]), //VTCʱ��������de��Ч��������
 .I_vtc_vs(I_vtc_vs),      //VTCʱ��������VSͬ���ź�����
 .I_vtc_vcnt(vcnt),        //vtc������ƫ�ƣ���Ҫ���з������ݽ��е���
 .O_pixel_en(wave1_pixel_en), //������ʹ��
 .single_flag(single_flag),
 .trigger_line(trigger_line),
 .trigger_edge(trigger_edge)//0�����أ�1�½���
 );
 /*
 //���λ���2���Լ����λ������ص����ʹ��
 uiwave_buf uiwave2_buf_inst
 (
 .I_wave_clk(I_wave2_clk),   //д��������ʱ�ӣ���ADC�ɼ�ʱ��ͬ��
 .I_wave_data(I_wave2_data), //д����
 .I_wave_data_de(I_wave2_data_de),//д������Ч
 .I_vtc_clk(I_vtc_clk),           //VTCʱ������ʱ������
 .I_vtc_rstn(I_vtc_rstn),         //VTCʱ��������λ 
 .I_vtc_de_r(vtc_de_r[0]),        //VTCʱ��������de��Ч��������
 .I_vtc_vs(I_vtc_vs),             //VTCʱ��������VSͬ���ź�����
 .I_vtc_vcnt(vcnt),               //vtc������ƫ�ƣ���Ҫ���з������ݽ��е���
 .O_pixel_en(wave2_pixel_en),      //������ʹ��
.single_flag(single_flag)
 );
 */
 endmodule