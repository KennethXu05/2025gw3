 module uiwave_buf
 (
 input         I_wave_clk,    //д��������ʱ�ӣ���ADC�ɼ�ʱ��ͬ��
 input  [7 :0] I_wave_data,   //д����
 input         I_wave_data_de,//д������Ч
 input         I_vtc_clk,     //VTCʱ������ʱ������
 input         I_vtc_rstn,    //VTCʱ��������λ 
 input         I_vtc_vs,      //VTCʱ��������VSͬ���ź�����
 input         I_vtc_de_r,    //VTCʱ��������de��Ч��������
 input  [7 :0] I_vtc_vcnt,    //vtc������ƫ�ƣ���Ҫ���з������ݽ��е���
 output        O_pixel_en,     //������ʹ��
 input         single_flag,
 input  [7:0 ] trigger_line,
 input         trigger_edge//0�����أ�1�½���

 );
 
 //BRAM ��˫��BRAM
 reg  [9 :0] addra = 0;  //BRAM ͨ��A��ַ     
 //reg         ena   = 0;  //BRAM ͨ��Aʹ�� 
 reg         wea   = 0;  //BRAM ͨ��Aдʹ��
 reg  [9 :0] addrb = 0;  //BRAM ͨ��B��ַ
 reg         enb   = 0;  //BRAM ͨ��B��ʹ��
 reg  [0 :0] WR_S,RD_S;  //д״̬������״̬��
 reg         buf_flag;//buf_flag����ƹ�ҵ�ַ�����л�
 reg         addr0_en;//��������д��һ��������Ե�ַ0
 
 wire [7 :0] wave_data;//д�������ݵ�BRAM
 reg  [3 :0] async_vtc_vs =0; //ͬ���ź�
 reg        trigger_select;
 always @(posedge I_wave_clk)begin //���첽I_vtc_vs����
     async_vtc_vs <= {async_vtc_vs[2:0],I_vtc_vs};
 end
 reg wave_data_de;
 reg [7:0]r_I_wave_data;
 always @(posedge I_wave_clk or negedge I_vtc_rstn) begin
    if(I_vtc_rstn == 1'b0)
      r_I_wave_data<=0;
    else
      r_I_wave_data<=I_wave_data;
 end

 wire trigger_flag;
 /*wire I_wave_data_around_min;
 wire I_wave_data_around_max;
 assign I_wave_data_around_max=(I_wave_data>=250)?255:I_wave_data+5;
 assign I_wave_data_around_min=(I_wave_data<=6)?1:I_wave_data-5; */
 assign trigger_flag=(trigger_line==I_wave_data)&&(((trigger_edge==0&&(r_I_wave_data<I_wave_data))||(trigger_edge==1)&&(r_I_wave_data>I_wave_data))?1'b1:1'b0);
 always @(posedge I_wave_clk or negedge I_vtc_rstn) begin
    if(I_vtc_rstn == 1'b0)begin
            wave_data_de<=0;
    end
    else if((WR_S==0)&&trigger_flag)begin
            wave_data_de<=I_wave_data_de;
    end
    else if(WR_S==1)begin
            wave_data_de<=0;
    end
    else
      wave_data_de<=wave_data_de;
 end
 //���Ʋ������ݵ�ʹ�ܣ�����ԭ��:
 //��ƥ�䵽�洢��ADC���ݺ�����ɨ���Y����ֵһ�¾������ÿ��X���귽�����1�����ε�

 assign   O_pixel_en  = I_vtc_de_r&(I_vtc_vcnt[7:0] == wave_data[7:0]);
 
 reg [21:0]trigger_cnt;
 always @(posedge I_wave_clk or negedge I_vtc_rstn) begin
    if(I_vtc_rstn == 1'b0)
      trigger_cnt<=0;
    else if((WR_S==0)&&trigger_flag)
      trigger_cnt<=0;
    else if(trigger_cnt>=22'd3_333_332)
      trigger_cnt<=trigger_cnt;
    else
      trigger_cnt<=trigger_cnt+1;
 end
 always @(posedge I_wave_clk or negedge I_vtc_rstn) begin
    if(I_vtc_rstn == 1'b0)begin
      trigger_select<=0;
    end
    else if((WR_S==0)&&trigger_flag)begin
      trigger_select<=1;
    end
    else if(trigger_cnt>=22'd3_333_332)begin
      trigger_select<=0;
    end
    else
      trigger_select<=trigger_select;
 end
 wire r_wave_data_de;
 assign r_wave_data_de=(trigger_select)?wave_data_de:I_wave_data_de;
 //дBRAM ״̬��
 always @(posedge I_wave_clk or negedge I_vtc_rstn)begin
     if(I_vtc_rstn == 1'b0)begin //��λ�������мĴ���
        addra      <= 10'd0;
        addr0_en   <= 1'b1;
        wea        <= 1'b0; 
        buf_flag   <= 1'b0;
        WR_S       <= 1'd0;
     end
     else begin
         case(WR_S) //д״̬��
         0:begin 
               if(r_wave_data_de)begin //��Ч�������ݵ�
                if(addra == 749)begin //1024������д��
                  wea      <= 1'b0; //ֹͣд
                  addra    <= 0;    //��Ե�ַ����0
                  addr0_en <= 1'b1;
                  WR_S     <= 1'd1;//����״̬��1
                end
                else begin //д��1024������
                  wea      <= 1'b1; //дʹ��
                  addr0_en <= 1'b0;
                  addra    <= (addr0_en == 1'b0) ? (addra + 1'b1) : 0;//��Ե�ַ����
                end
             end
             else begin
               wea <= 1'b0;
             end
         end
         1:begin //�ȴ�VTCʱ��ͬ��
             if(single_flag)begin
                buf_flag<=buf_flag;
                if(async_vtc_vs[3:2] == 2'b10)begin//������ͬ����׼����һ��д
                WR_S     <= 1'd0; //�ص�״̬0
             end
             end
             else if(async_vtc_vs[3:2] == 2'b10)begin//������ͬ����׼����һ��д
                WR_S     <= 1'd0; //�ص�״̬0
                buf_flag <= ~buf_flag;//ƹ�ҵ�ַ�л�
             end
         end
         default:WR_S   <= 2'd0;
         endcase
      end
 end
 
 //��BRAM ״̬��
 always @(posedge I_vtc_clk or negedge I_vtc_rstn)begin
     if(I_vtc_rstn == 1'b0)begin//��λ�������мĴ���
        addrb   <= 10'd0;
        RD_S    <= 1'd0;
     end
     else begin
         case(RD_S)
         0:begin
             if(I_vtc_de_r)begin //I_vtc_de_r��������Ч��������
                if(addrb == 749)begin //1024�����ݶ���
                  addrb <= 0;    //��Ե�ַ����0
                  RD_S  <= 1'd1; //����״̬1
                end
                else //ûһ������ɨ�����е�ADC����
                  addrb   <= addrb + 1'b1;//��Ե�ַ����
             end
         end
         1:begin
             if(I_vtc_de_r == 0) //�ȴ�de��Ϊ0
                 RD_S <= 0; //�ص�״̬0����ɨ��
                 
         end
         default:RD_S   <= 1'd0;
         endcase
      end
 end   
 wave_ram buf_inst(
        .dout(wave_data), //output [7:0] dout
        .clka(I_wave_clk), //input clka
        .cea(wea), //input cea
        .clkb(I_vtc_clk), //input clkb
        .ceb(1'b1), //input ceb
        .oce(1'b1), //input oce
        .reset(!I_vtc_rstn), //input reset
        .ada({buf_flag,addra}), //input [9:0] ada
        .din(I_wave_data), //input [7:0] din
        .adb({~buf_flag,addrb}) //input [9:0] adb
    );/*
 wave_ram buf_inst( 
 .dina(I_wave_data), //д�벨������
 .addra({buf_flag,addra}), //д��ַ������addra����Ե�ַ��buf_flag�ǵ�ַ��λ�����ڶ�д��ƹ���л�
 .wea(wea), //дʹ��
 .clka(I_wave_clk),//дʱ��
 .doutb(wave_data), //�����Ĳ�������
 .addrb({~buf_flag,addrb}), //д��ַ������addrb����Ե�ַ��buf_flag�ǵ�ַ��λ�����ڶ�д��ƹ���л�
 .clkb(I_vtc_clk)//��ʱ��
 );*/
 endmodule