//Copyright (C)2014-2025 Gowin Semiconductor Corporation.
//All rights reserved.
//File Title: IP file
//Tool Version: V1.9.12 (64-bit)
//Part Number: GW5AT-LV138PG484AC1/I0
//Device: GW5AT-138
//Device Version: B
//Created Time: Thu Oct  9 14:53:57 2025

module tri_pROM (dout, clk, oce, ce, reset, ad);

output [7:0] dout;
input clk;
input oce;
input ce;
input reset;
input [10:0] ad;

wire [23:0] prom_inst_0_dout_w;
wire gw_gnd;

assign gw_gnd = 1'b0;

pROM prom_inst_0 (
    .DO({prom_inst_0_dout_w[23:0],dout[7:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .AD({ad[10:0],gw_gnd,gw_gnd,gw_gnd})
);

defparam prom_inst_0.READ_MODE = 1'b0;
defparam prom_inst_0.BIT_WIDTH = 8;
defparam prom_inst_0.RESET_MODE = "SYNC";
defparam prom_inst_0.INIT_RAM_00 = 256'h0D0C0C0B0B0B0A0A090909080807070706060505040404030302020201010000;
defparam prom_inst_0.INIT_RAM_01 = 256'h1A191919181817171616161515141414131312121211111010100F0F0E0E0D0D;
defparam prom_inst_0.INIT_RAM_02 = 256'h2726262625252424242323222222212120201F1F1F1E1E1D1D1D1C1C1B1B1B1A;
defparam prom_inst_0.INIT_RAM_03 = 256'h34333333323231313130302F2F2F2E2E2D2D2D2C2C2B2B2B2A2A292928282827;
defparam prom_inst_0.INIT_RAM_04 = 256'h414140403F3F3F3E3E3D3D3C3C3C3B3B3A3A3A39393838383737363636353534;
defparam prom_inst_0.INIT_RAM_05 = 256'h4E4E4D4D4C4C4C4B4B4A4A4A4949484848474746464545454444434343424241;
defparam prom_inst_0.INIT_RAM_06 = 256'h5B5B5A5A595959585857575756565555555454535353525251515150504F4F4E;
defparam prom_inst_0.INIT_RAM_07 = 256'h686867676766666565656464636362626261616060605F5F5E5E5E5D5D5C5C5C;
defparam prom_inst_0.INIT_RAM_08 = 256'h7575747474737372727271717070706F6F6E6E6E6D6D6C6C6B6B6B6A6A696969;
defparam prom_inst_0.INIT_RAM_09 = 256'h82828281818080807F7F7E7E7D7D7D7C7C7B7B7B7A7A79797978787777777676;
defparam prom_inst_0.INIT_RAM_0A = 256'h8F8F8F8E8E8D8D8D8C8C8B8B8B8A8A8989888888878786868685858484848383;
defparam prom_inst_0.INIT_RAM_0B = 256'h9D9C9C9B9B9A9A9A999998989897979696969595949494939392929191919090;
defparam prom_inst_0.INIT_RAM_0C = 256'hAAA9A9A8A8A8A7A7A6A6A6A5A5A4A4A3A3A3A2A2A1A1A1A0A09F9F9F9E9E9D9D;
defparam prom_inst_0.INIT_RAM_0D = 256'hB7B6B6B5B5B5B4B4B3B3B3B2B2B1B1B1B0B0AFAFAEAEAEADADACACACABABAAAA;
defparam prom_inst_0.INIT_RAM_0E = 256'hC4C3C3C3C2C2C1C1C0C0C0BFBFBEBEBEBDBDBCBCBCBBBBBABABAB9B9B8B8B7B7;
defparam prom_inst_0.INIT_RAM_0F = 256'hD1D0D0D0CFCFCECECECDCDCCCCCCCBCBCACAC9C9C9C8C8C7C7C7C6C6C5C5C5C4;
defparam prom_inst_0.INIT_RAM_10 = 256'hDEDDDDDDDCDCDBDBDBDADAD9D9D9D8D8D7D7D7D6D6D5D5D5D4D4D3D3D2D2D2D1;
defparam prom_inst_0.INIT_RAM_11 = 256'hEBEBEAEAE9E9E9E8E8E7E7E6E6E6E5E5E4E4E4E3E3E2E2E2E1E1E0E0E0DFDFDE;
defparam prom_inst_0.INIT_RAM_12 = 256'hF8F8F7F7F6F6F6F5F5F4F4F4F3F3F2F2F2F1F1F0F0EFEFEFEEEEEDEDEDECECEB;
defparam prom_inst_0.INIT_RAM_13 = 256'hF9FAFAFBFBFBFCFCFDFDFDFEFEFFFFFFFFFEFEFDFDFDFCFCFBFBFBFAFAF9F9F8;
defparam prom_inst_0.INIT_RAM_14 = 256'hECEDEDEDEEEEEFEFEFF0F0F1F1F2F2F2F3F3F4F4F4F5F5F6F6F6F7F7F8F8F8F9;
defparam prom_inst_0.INIT_RAM_15 = 256'hDFE0E0E0E1E1E2E2E2E3E3E4E4E4E5E5E6E6E6E7E7E8E8E9E9E9EAEAEBEBEBEC;
defparam prom_inst_0.INIT_RAM_16 = 256'hD2D2D3D3D4D4D5D5D5D6D6D7D7D7D8D8D9D9D9DADADBDBDBDCDCDDDDDDDEDEDF;
defparam prom_inst_0.INIT_RAM_17 = 256'hC5C5C6C6C7C7C7C8C8C9C9C9CACACBCBCCCCCCCDCDCECECECFCFD0D0D0D1D1D2;
defparam prom_inst_0.INIT_RAM_18 = 256'hB8B8B9B9BABABABBBBBCBCBCBDBDBEBEBEBFBFC0C0C0C1C1C2C2C3C3C3C4C4C5;
defparam prom_inst_0.INIT_RAM_19 = 256'hABABACACACADADAEAEAEAFAFB0B0B1B1B1B2B2B3B3B3B4B4B5B5B5B6B6B7B7B7;
defparam prom_inst_0.INIT_RAM_1A = 256'h9E9E9F9F9FA0A0A1A1A1A2A2A3A3A3A4A4A5A5A6A6A6A7A7A8A8A8A9A9AAAAAA;
defparam prom_inst_0.INIT_RAM_1B = 256'h919191929293939494949595969696979798989899999A9A9A9B9B9C9C9D9D9D;
defparam prom_inst_0.INIT_RAM_1C = 256'h8484848585868686878788888889898A8A8B8B8B8C8C8D8D8D8E8E8F8F8F9090;
defparam prom_inst_0.INIT_RAM_1D = 256'h77777778787979797A7A7B7B7B7C7C7D7D7D7E7E7F7F80808081818282828383;
defparam prom_inst_0.INIT_RAM_1E = 256'h696A6A6B6B6B6C6C6D6D6E6E6E6F6F7070707171727272737374747475757676;
defparam prom_inst_0.INIT_RAM_1F = 256'h5C5D5D5E5E5E5F5F606060616162626263636464656565666667676768686969;
defparam prom_inst_0.INIT_RAM_20 = 256'h4F505051515152525353535454555555565657575758585959595A5A5B5B5C5C;
defparam prom_inst_0.INIT_RAM_21 = 256'h4243434344444545454646474748484849494A4A4A4B4B4C4C4C4D4D4E4E4E4F;
defparam prom_inst_0.INIT_RAM_22 = 256'h35363636373738383839393A3A3A3B3B3C3C3C3D3D3E3E3F3F3F404041414142;
defparam prom_inst_0.INIT_RAM_23 = 256'h282829292A2A2B2B2B2C2C2D2D2D2E2E2F2F2F30303131313232333333343435;
defparam prom_inst_0.INIT_RAM_24 = 256'h1B1B1C1C1D1D1D1E1E1F1F1F2020212122222223232424242525262626272728;
defparam prom_inst_0.INIT_RAM_25 = 256'h0E0E0F0F101010111112121213131414141515161616171718181919191A1A1B;
defparam prom_inst_0.INIT_RAM_26 = 256'h010102020203030404040505060607070708080909090A0A0B0B0B0C0C0D0D0D;
defparam prom_inst_0.INIT_RAM_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;

endmodule //tri_pROM
