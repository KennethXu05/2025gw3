//Copyright (C)2014-2025 Gowin Semiconductor Corporation.
//All rights reserved.
//File Title: IP file
//Tool Version: V1.9.12 (64-bit)
//Part Number: GW5AT-LV138PG484AC1/I0
//Device: GW5AT-138
//Device Version: B
//Created Time: Fri Oct  3 12:06:57 2025

module Gowin_pROM_spwm_sin (dout, clk, oce, ce, reset, ad);

output [9:0] dout;
input clk;
input oce;
input ce;
input reset;
input [9:0] ad;

wire [21:0] prom_inst_0_dout_w;
wire gw_gnd;

assign gw_gnd = 1'b0;

pROM prom_inst_0 (
    .DO({prom_inst_0_dout_w[21:0],dout[9:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .AD({ad[9:0],gw_gnd,gw_gnd,gw_gnd,gw_gnd})
);

defparam prom_inst_0.READ_MODE = 1'b0;
defparam prom_inst_0.BIT_WIDTH = 16;
defparam prom_inst_0.RESET_MODE = "SYNC";
defparam prom_inst_0.INIT_RAM_00 = 256'h022F022C022902250222021F021C021902150212020F020C02090205020201FF;
defparam prom_inst_0.INIT_RAM_01 = 256'h0262025F025C025802550252024F024C024902450242023F023C023902350232;
defparam prom_inst_0.INIT_RAM_02 = 256'h02940291028E028A028702840281027E027B027802750272026E026B02680265;
defparam prom_inst_0.INIT_RAM_03 = 256'h02C402C102BE02BB02B802B502B202AF02AC02A902A602A302A0029D029A0297;
defparam prom_inst_0.INIT_RAM_04 = 256'h02F202F002ED02EA02E702E402E102DE02DB02D902D602D302D002CD02CA02C7;
defparam prom_inst_0.INIT_RAM_05 = 256'h031E031C0319031603140311030E030B030903060303030002FE02FB02F802F5;
defparam prom_inst_0.INIT_RAM_06 = 256'h0347034503420340033D033B0338033603330331032E032B0329032603240321;
defparam prom_inst_0.INIT_RAM_07 = 256'h036D036B0368036603640361035F035D035A0358035603530351034F034C034A;
defparam prom_inst_0.INIT_RAM_08 = 256'h038F038D038B03890387038503830380037E037C037A0378037603740371036F;
defparam prom_inst_0.INIT_RAM_09 = 256'h03AD03AB03A903A703A603A403A203A0039E039C039B03990397039503930391;
defparam prom_inst_0.INIT_RAM_0A = 256'h03C603C503C303C203C003BF03BD03BC03BA03B803B703B503B403B203B003AE;
defparam prom_inst_0.INIT_RAM_0B = 256'h03DB03DA03D903D803D603D503D403D303D103D003CF03CD03CC03CB03C903C8;
defparam prom_inst_0.INIT_RAM_0C = 256'h03EB03EB03EA03E903E803E703E603E503E403E303E203E103E003DF03DE03DC;
defparam prom_inst_0.INIT_RAM_0D = 256'h03F703F603F603F503F403F403F303F203F203F103F003F003EF03EE03ED03EC;
defparam prom_inst_0.INIT_RAM_0E = 256'h03FD03FD03FC03FC03FC03FB03FB03FB03FA03FA03FA03F903F903F803F803F7;
defparam prom_inst_0.INIT_RAM_0F = 256'h03FE03FE03FE03FE03FE03FE03FE03FE03FE03FE03FE03FE03FE03FD03FD03FD;
defparam prom_inst_0.INIT_RAM_10 = 256'h03FA03FA03FA03FB03FB03FB03FC03FC03FC03FD03FD03FD03FD03FD03FE03FE;
defparam prom_inst_0.INIT_RAM_11 = 256'h03F003F103F203F203F303F403F403F503F603F603F703F703F803F803F903F9;
defparam prom_inst_0.INIT_RAM_12 = 256'h03E203E303E403E503E603E703E803E903EA03EB03EB03EC03ED03EE03EF03F0;
defparam prom_inst_0.INIT_RAM_13 = 256'h03CF03D003D103D303D403D503D603D803D903DA03DB03DC03DE03DF03E003E1;
defparam prom_inst_0.INIT_RAM_14 = 256'h03B703B803BA03BC03BD03BF03C003C203C303C503C603C803C903CB03CC03CD;
defparam prom_inst_0.INIT_RAM_15 = 256'h039B039C039E03A003A203A403A603A703A903AB03AD03AE03B003B203B403B5;
defparam prom_inst_0.INIT_RAM_16 = 256'h037A037C037E03800383038503870389038B038D038F03910393039503970399;
defparam prom_inst_0.INIT_RAM_17 = 256'h03560358035A035D035F0361036403660368036B036D036F0371037403760378;
defparam prom_inst_0.INIT_RAM_18 = 256'h032E0331033303360338033B033D0340034203450347034A034C034F03510353;
defparam prom_inst_0.INIT_RAM_19 = 256'h030303060309030B030E0311031403160319031C031E0321032403260329032B;
defparam prom_inst_0.INIT_RAM_1A = 256'h02D602D902DB02DE02E102E402E702EA02ED02F002F202F502F802FB02FE0300;
defparam prom_inst_0.INIT_RAM_1B = 256'h02A602A902AC02AF02B202B502B802BB02BE02C102C402C702CA02CD02D002D3;
defparam prom_inst_0.INIT_RAM_1C = 256'h02750278027B027E028102840287028A028E029102940297029A029D02A002A3;
defparam prom_inst_0.INIT_RAM_1D = 256'h024202450249024C024F025202550258025C025F026202650268026B026E0272;
defparam prom_inst_0.INIT_RAM_1E = 256'h020F021202150219021C021F022202250229022C022F023202350239023C023F;
defparam prom_inst_0.INIT_RAM_1F = 256'h01DC01DF01E201E501E901EC01EF01F201F501F901FC01FF020202050209020C;
defparam prom_inst_0.INIT_RAM_20 = 256'h01A901AC01AF01B201B501B901BC01BF01C201C501C901CC01CF01D201D501D9;
defparam prom_inst_0.INIT_RAM_21 = 256'h0177017A017D0180018301860189018C0190019301960199019C019F01A201A6;
defparam prom_inst_0.INIT_RAM_22 = 256'h01460149014C014F015201550158015B015E016101640167016A016D01700174;
defparam prom_inst_0.INIT_RAM_23 = 256'h0117011A011D0120012301250128012B012E013101340137013A013D01400143;
defparam prom_inst_0.INIT_RAM_24 = 256'h00EA00ED00F000F300F500F800FB00FE0100010301060109010C010E01110114;
defparam prom_inst_0.INIT_RAM_25 = 256'h00C100C300C600C800CB00CD00D000D300D500D800DA00DD00E000E200E500E8;
defparam prom_inst_0.INIT_RAM_26 = 256'h009A009D009F00A100A400A600A800AB00AD00AF00B200B400B700B900BC00BE;
defparam prom_inst_0.INIT_RAM_27 = 256'h00770079007B007E00800082008400860088008A008D008F0091009300960098;
defparam prom_inst_0.INIT_RAM_28 = 256'h0058005A005C005E006000620063006500670069006B006D006F007100730075;
defparam prom_inst_0.INIT_RAM_29 = 256'h003E003F004100420044004600470049004A004C004E00500051005300550057;
defparam prom_inst_0.INIT_RAM_2A = 256'h00280029002A002B002D002E002F0031003200330035003600380039003B003C;
defparam prom_inst_0.INIT_RAM_2B = 256'h0016001700180019001A001B001C001D001E001F002000220023002400250026;
defparam prom_inst_0.INIT_RAM_2C = 256'h000A000A000B000C000C000D000E000E000F0010001100120013001300140015;
defparam prom_inst_0.INIT_RAM_2D = 256'h0002000300030003000400040004000500050006000600070007000800080009;
defparam prom_inst_0.INIT_RAM_2E = 256'h0000000000000000000000000000000000000001000100010001000100020002;
defparam prom_inst_0.INIT_RAM_2F = 256'h0003000300020002000200010001000100010001000000000000000000000000;
defparam prom_inst_0.INIT_RAM_30 = 256'h000B000A000A0009000800080007000700060006000500050004000400040003;
defparam prom_inst_0.INIT_RAM_31 = 256'h0018001700160015001400130013001200110010000F000E000E000D000C000C;
defparam prom_inst_0.INIT_RAM_32 = 256'h002A00290028002600250024002300220020001F001E001D001C001B001A0019;
defparam prom_inst_0.INIT_RAM_33 = 256'h0041003F003E003C003B0039003800360035003300320031002F002E002D002B;
defparam prom_inst_0.INIT_RAM_34 = 256'h005C005A005800570055005300510050004E004C004A00490047004600440042;
defparam prom_inst_0.INIT_RAM_35 = 256'h007B00790077007500730071006F006D006B006900670065006300620060005E;
defparam prom_inst_0.INIT_RAM_36 = 256'h009F009D009A0098009600930091008F008D008A00880086008400820080007E;
defparam prom_inst_0.INIT_RAM_37 = 256'h00C600C300C100BE00BC00B900B700B400B200AF00AD00AB00A800A600A400A1;
defparam prom_inst_0.INIT_RAM_38 = 256'h00F000ED00EA00E800E500E200E000DD00DA00D800D500D300D000CD00CB00C8;
defparam prom_inst_0.INIT_RAM_39 = 256'h011D011A011701140111010E010C010901060103010000FE00FB00F800F500F3;
defparam prom_inst_0.INIT_RAM_3A = 256'h014C0149014601430140013D013A013701340131012E012B0128012501230120;
defparam prom_inst_0.INIT_RAM_3B = 256'h017D017A017701740170016D016A016701640161015E015B015801550152014F;
defparam prom_inst_0.INIT_RAM_3C = 256'h01AF01AC01A901A601A2019F019C0199019601930190018C0189018601830180;
defparam prom_inst_0.INIT_RAM_3D = 256'h01E201DF01DC01D901D501D201CF01CC01C901C501C201BF01BC01B901B501B2;
defparam prom_inst_0.INIT_RAM_3E = 256'h0000000000000000000000000000000001FC01F901F501F201EF01EC01E901E5;

endmodule //Gowin_pROM_spwm_sin
