//Copyright (C)2014-2025 Gowin Semiconductor Corporation.
//All rights reserved.
//File Title: IP file
//Tool Version: V1.9.12 (64-bit)
//Part Number: GW5AT-LV138PG484AC1/I0
//Device: GW5AT-138
//Device Version: B
//Created Time: Thu Oct  9 14:48:05 2025

module sin_pROM (dout, clk, oce, ce, reset, ad);

output [7:0] dout;
input clk;
input oce;
input ce;
input reset;
input [10:0] ad;

wire [23:0] prom_inst_0_dout_w;
wire gw_gnd;

assign gw_gnd = 1'b0;

pROM prom_inst_0 (
    .DO({prom_inst_0_dout_w[23:0],dout[7:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .AD({ad[10:0],gw_gnd,gw_gnd,gw_gnd})
);

defparam prom_inst_0.READ_MODE = 1'b0;
defparam prom_inst_0.BIT_WIDTH = 8;
defparam prom_inst_0.RESET_MODE = "SYNC";
defparam prom_inst_0.INIT_RAM_00 = 256'h9392919190908F8E8E8D8C8C8B8A8A898988878786858584838382828180807F;
defparam prom_inst_0.INIT_RAM_01 = 256'hA7A6A5A5A4A4A3A2A2A1A0A09F9F9E9D9D9C9B9B9A9A99989897969695959493;
defparam prom_inst_0.INIT_RAM_02 = 256'hB9B9B8B8B7B7B6B5B5B4B4B3B2B2B1B1B0B0AFAEAEADADACABABAAAAA9A8A8A7;
defparam prom_inst_0.INIT_RAM_03 = 256'hCBCACAC9C9C8C8C7C7C6C5C5C4C4C3C3C2C2C1C1C0C0BFBEBEBDBDBCBCBBBABA;
defparam prom_inst_0.INIT_RAM_04 = 256'hDADAD9D9D8D8D7D7D6D6D5D5D5D4D4D3D3D2D2D1D1D0D0CFCFCECECDCDCCCCCB;
defparam prom_inst_0.INIT_RAM_05 = 256'hE7E7E6E6E6E5E5E4E4E4E3E3E2E2E2E1E1E0E0E0DFDFDEDEDEDDDDDCDCDBDBDA;
defparam prom_inst_0.INIT_RAM_06 = 256'hF1F1F1F1F0F0F0EFEFEFEEEEEEEEEDEDEDECECECEBEBEBEAEAEAE9E9E8E8E8E7;
defparam prom_inst_0.INIT_RAM_07 = 256'hF9F9F8F8F8F8F8F7F7F7F7F7F6F6F6F6F5F5F5F5F4F4F4F4F3F3F3F3F2F2F2F2;
defparam prom_inst_0.INIT_RAM_08 = 256'hFDFDFDFDFDFDFCFCFCFCFCFCFCFCFCFBFBFBFBFBFBFBFAFAFAFAFAFAF9F9F9F9;
defparam prom_inst_0.INIT_RAM_09 = 256'hFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFEFDFDFDFDFDFDFD;
defparam prom_inst_0.INIT_RAM_0A = 256'hFCFCFCFCFCFCFCFCFDFDFDFDFDFDFDFDFDFDFDFDFDFEFEFEFEFEFEFEFEFEFEFE;
defparam prom_inst_0.INIT_RAM_0B = 256'hF6F6F7F7F7F7F7F8F8F8F8F8F9F9F9F9F9F9FAFAFAFAFAFAFBFBFBFBFBFBFBFC;
defparam prom_inst_0.INIT_RAM_0C = 256'hEEEEEEEEEFEFEFF0F0F0F1F1F1F1F2F2F2F2F3F3F3F3F4F4F4F4F5F5F5F5F6F6;
defparam prom_inst_0.INIT_RAM_0D = 256'hE2E2E3E3E4E4E4E5E5E6E6E6E7E7E7E8E8E8E9E9EAEAEAEBEBEBECECECEDEDED;
defparam prom_inst_0.INIT_RAM_0E = 256'hD4D5D5D5D6D6D7D7D8D8D9D9DADADADBDBDCDCDDDDDEDEDEDFDFE0E0E0E1E1E2;
defparam prom_inst_0.INIT_RAM_0F = 256'hC4C4C5C5C6C7C7C8C8C9C9CACACBCBCCCCCDCDCECECFCFD0D0D1D1D2D2D3D3D4;
defparam prom_inst_0.INIT_RAM_10 = 256'hB2B2B3B4B4B5B5B6B7B7B8B8B9B9BABABBBCBCBDBDBEBEBFC0C0C1C1C2C2C3C3;
defparam prom_inst_0.INIT_RAM_11 = 256'h9F9FA0A0A1A2A2A3A4A4A5A5A6A7A7A8A8A9AAAAABABACADADAEAEAFB0B0B1B1;
defparam prom_inst_0.INIT_RAM_12 = 256'h8A8B8C8C8D8E8E8F909091919293939495959696979898999A9A9B9B9C9D9D9E;
defparam prom_inst_0.INIT_RAM_13 = 256'h7677777879797A7B7B7C7C7D7E7E7F808081828283838485858687878889898A;
defparam prom_inst_0.INIT_RAM_14 = 256'h626363646465666667686869696A6B6B6C6D6D6E6E6F70707172727374747575;
defparam prom_inst_0.INIT_RAM_15 = 256'h4E4F50505151525353545455565657575859595A5A5B5C5C5D5E5E5F5F606161;
defparam prom_inst_0.INIT_RAM_16 = 256'h3C3D3D3E3E3F4040414142424344444545464647474849494A4A4B4C4C4D4D4E;
defparam prom_inst_0.INIT_RAM_17 = 256'h2C2C2D2D2E2E2F2F303031313232333334343535363637373839393A3A3B3B3C;
defparam prom_inst_0.INIT_RAM_18 = 256'h1E1E1E1F1F20202021212222232324242425252626272728282929292A2A2B2B;
defparam prom_inst_0.INIT_RAM_19 = 256'h121212131313141414151516161617171718181819191A1A1A1B1B1C1C1C1D1D;
defparam prom_inst_0.INIT_RAM_1A = 256'h0909090A0A0A0A0B0B0B0B0C0C0C0C0D0D0D0D0E0E0E0F0F0F10101010111111;
defparam prom_inst_0.INIT_RAM_1B = 256'h0303030303040404040404050505050505060606060607070707070808080809;
defparam prom_inst_0.INIT_RAM_1C = 256'h0000000000000000010101010101010101010101010202020202020202020303;
defparam prom_inst_0.INIT_RAM_1D = 256'h0101010100000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_1E = 256'h0504040404040403030303030303020202020202020202010101010101010101;
defparam prom_inst_0.INIT_RAM_1F = 256'h0C0B0B0B0B0A0A0A0A0909090908080808070707070706060606060505050505;
defparam prom_inst_0.INIT_RAM_20 = 256'h161515141414131313121212111111101010100F0F0F0E0E0E0D0D0D0D0C0C0C;
defparam prom_inst_0.INIT_RAM_21 = 256'h222221212020201F1F1E1E1E1D1D1C1C1C1B1B1A1A1A19191818181717171616;
defparam prom_inst_0.INIT_RAM_22 = 256'h313130302F2F2E2E2D2D2C2C2B2B2A2A29292928282727262625252424242323;
defparam prom_inst_0.INIT_RAM_23 = 256'h4242414140403F3E3E3D3D3C3C3B3B3A3A393938373736363535343433333232;
defparam prom_inst_0.INIT_RAM_24 = 256'h555454535352515150504F4E4E4D4D4C4C4B4A4A494948474746464545444443;
defparam prom_inst_0.INIT_RAM_25 = 256'h6968686766666564646363626161605F5F5E5E5D5C5C5B5A5A59595857575656;
defparam prom_inst_0.INIT_RAM_26 = 256'h7D7C7C7B7B7A797978777776757574747372727170706F6E6E6D6D6C6B6B6A69;
defparam prom_inst_0.INIT_RAM_27 = 256'h0000000000000000000000000000000000000000000000000000000000007E7E;

endmodule //sin_pROM
