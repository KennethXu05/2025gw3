//Copyright (C)2014-2025 Gowin Semiconductor Corporation.
//All rights reserved.
//File Title: IP file
//Tool Version: V1.9.12 (64-bit)
//Part Number: GW5AT-LV138PG484AC1/I0
//Device: GW5AT-138
//Device Version: B
//Created Time: Thu Oct  9 14:56:38 2025

module saw_pROM (dout, clk, oce, ce, reset, ad);

output [7:0] dout;
input clk;
input oce;
input ce;
input reset;
input [10:0] ad;

wire [23:0] prom_inst_0_dout_w;
wire gw_gnd;

assign gw_gnd = 1'b0;

pROM prom_inst_0 (
    .DO({prom_inst_0_dout_w[23:0],dout[7:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .AD({ad[10:0],gw_gnd,gw_gnd,gw_gnd})
);

defparam prom_inst_0.READ_MODE = 1'b0;
defparam prom_inst_0.BIT_WIDTH = 8;
defparam prom_inst_0.RESET_MODE = "SYNC";
defparam prom_inst_0.INIT_RAM_00 = 256'h0808070707070606060605050505040404040303030302020202010101010000;
defparam prom_inst_0.INIT_RAM_01 = 256'h1010100F0F0F0F0E0E0E0E0D0D0D0D0C0C0C0B0B0B0B0A0A0A0A090909090808;
defparam prom_inst_0.INIT_RAM_02 = 256'h1818181717171716161616151515151414141413131313121212121111111110;
defparam prom_inst_0.INIT_RAM_03 = 256'h202020201F1F1F1F1E1E1E1E1D1D1D1D1C1C1C1C1B1B1B1B1A1A1A1A19191919;
defparam prom_inst_0.INIT_RAM_04 = 256'h2928282828272727272626262625252525242424232323232222222221212121;
defparam prom_inst_0.INIT_RAM_05 = 256'h31303030302F2F2F2F2E2E2E2E2D2D2D2D2C2C2C2C2B2B2B2B2A2A2A2A292929;
defparam prom_inst_0.INIT_RAM_06 = 256'h3939383838383737373736363636353535353434343433333333323232323131;
defparam prom_inst_0.INIT_RAM_07 = 256'h414141404040403F3F3F3F3E3E3E3E3D3D3D3C3C3C3C3B3B3B3B3A3A3A3A3939;
defparam prom_inst_0.INIT_RAM_08 = 256'h4949494848484847474747464646464545454544444444434343434242424241;
defparam prom_inst_0.INIT_RAM_09 = 256'h51515151505050504F4F4F4F4E4E4E4E4D4D4D4D4C4C4C4C4B4B4B4B4A4A4A4A;
defparam prom_inst_0.INIT_RAM_0A = 256'h5A59595959585858585757575756565656555555545454545353535352525252;
defparam prom_inst_0.INIT_RAM_0B = 256'h6262616161606060605F5F5F5F5E5E5E5E5D5D5D5D5C5C5C5C5B5B5B5B5A5A5A;
defparam prom_inst_0.INIT_RAM_0C = 256'h6A6A696969696868686867676767666666666565656564646464636363636262;
defparam prom_inst_0.INIT_RAM_0D = 256'h72727271717171707070706F6F6F6F6E6E6E6E6D6D6D6C6C6C6C6B6B6B6B6A6A;
defparam prom_inst_0.INIT_RAM_0E = 256'h7A7A7A7A79797978787878777777777676767675757575747474747373737372;
defparam prom_inst_0.INIT_RAM_0F = 256'h8282828281818181808080807F7F7F7F7E7E7E7E7D7D7D7D7C7C7C7C7B7B7B7B;
defparam prom_inst_0.INIT_RAM_10 = 256'h8B8A8A8A8A898989898888888887878787868686858585858484848483838383;
defparam prom_inst_0.INIT_RAM_11 = 256'h939392929291919191909090908F8F8F8F8E8E8E8E8D8D8D8D8C8C8C8C8B8B8B;
defparam prom_inst_0.INIT_RAM_12 = 256'h9B9B9A9A9A9A9999999998989898979797979696969695959595949494949393;
defparam prom_inst_0.INIT_RAM_13 = 256'hA3A3A3A2A2A2A2A1A1A1A1A0A0A0A09F9F9F9F9E9E9E9D9D9D9D9C9C9C9C9B9B;
defparam prom_inst_0.INIT_RAM_14 = 256'hABABABABAAAAAAA9A9A9A9A8A8A8A8A7A7A7A7A6A6A6A6A5A5A5A5A4A4A4A4A3;
defparam prom_inst_0.INIT_RAM_15 = 256'hB3B3B3B3B2B2B2B2B1B1B1B1B0B0B0B0AFAFAFAFAEAEAEAEADADADADACACACAC;
defparam prom_inst_0.INIT_RAM_16 = 256'hBCBBBBBBBBBABABABAB9B9B9B9B8B8B8B8B7B7B7B7B6B6B6B5B5B5B5B4B4B4B4;
defparam prom_inst_0.INIT_RAM_17 = 256'hC4C4C3C3C3C3C2C2C2C1C1C1C1C0C0C0C0BFBFBFBFBEBEBEBEBDBDBDBDBCBCBC;
defparam prom_inst_0.INIT_RAM_18 = 256'hCCCCCBCBCBCBCACACACAC9C9C9C9C8C8C8C8C7C7C7C7C6C6C6C6C5C5C5C5C4C4;
defparam prom_inst_0.INIT_RAM_19 = 256'hD4D4D4D3D3D3D3D2D2D2D2D1D1D1D1D0D0D0D0CFCFCFCFCECECECDCDCDCDCCCC;
defparam prom_inst_0.INIT_RAM_1A = 256'hDCDCDCDCDBDBDBDADADADAD9D9D9D9D8D8D8D8D7D7D7D7D6D6D6D6D5D5D5D5D4;
defparam prom_inst_0.INIT_RAM_1B = 256'hE4E4E4E4E3E3E3E3E2E2E2E2E1E1E1E1E0E0E0E0DFDFDFDFDEDEDEDEDDDDDDDD;
defparam prom_inst_0.INIT_RAM_1C = 256'hEDECECECECEBEBEBEBEAEAEAEAE9E9E9E9E8E8E8E8E7E7E7E6E6E6E6E5E5E5E5;
defparam prom_inst_0.INIT_RAM_1D = 256'hF5F5F4F4F4F4F3F3F3F2F2F2F2F1F1F1F1F0F0F0F0EFEFEFEFEEEEEEEEEDEDED;
defparam prom_inst_0.INIT_RAM_1E = 256'hFDFDFCFCFCFCFBFBFBFBFAFAFAFAF9F9F9F9F8F8F8F8F7F7F7F7F6F6F6F6F5F5;
defparam prom_inst_0.INIT_RAM_1F = 256'hE7E8E9EBECEDEEEFF0F1F2F3F4F5F6F7F8F9FAFBFCFDFEFFFFFFFEFEFEFEFDFD;
defparam prom_inst_0.INIT_RAM_20 = 256'hC7C8C9CACBCCCDCECFD0D1D2D3D4D5D6D7D8D9DADBDCDDDEDFE0E1E2E3E4E5E6;
defparam prom_inst_0.INIT_RAM_21 = 256'hA6A7A8A9AAABACADAEAFB0B1B2B3B4B5B6B7B8B9BABBBCBDBEC0C1C2C3C4C5C6;
defparam prom_inst_0.INIT_RAM_22 = 256'h85868788898A8B8C8D8E8F9091929394969798999A9B9C9D9E9FA0A1A2A3A4A5;
defparam prom_inst_0.INIT_RAM_23 = 256'h6465666768696B6C6D6E6F707172737475767778797A7B7C7D7E7F8081828384;
defparam prom_inst_0.INIT_RAM_24 = 256'h4445464748494A4B4C4D4E4F505152535455565758595A5B5C5D5E5F60616263;
defparam prom_inst_0.INIT_RAM_25 = 256'h232425262728292A2B2C2D2E2F303132333435363738393A3B3C3D3E3F414243;
defparam prom_inst_0.INIT_RAM_26 = 256'h02030405060708090A0B0C0D0E0F1011121314161718191A1B1C1D1E1F202122;
defparam prom_inst_0.INIT_RAM_27 = 256'h0000000000000000000000000000000000000000000000000000000000000001;

endmodule //saw_pROM
