module HDMI_PLL(
    clkin,
    init_clk,
    clkout0,
    clkout1,
    lock,
    reset
);


input clkin;
input init_clk;
output clkout0;
output clkout1;
output lock;
input reset;
wire [5:0] icpsel;
wire [2:0] lpfres;
wire pll_lock;
wire pll_rst;


    HDMI_PLL_MOD u_pll_HDMI(
        .clkout1(clkout1),
        .clkout0(clkout0),
        .lock(pll_lock),
        .clkin(clkin),
        .reset(pll_rst),
        .icpsel(icpsel),
        .lpfres(lpfres),
        .lpfcap(2'b00)
    );


    PLL_INIT_HDMI u_pll_init_HDMI(
        .CLKIN(init_clk),
        .I_RST(reset),
        .O_RST(pll_rst),
        .PLLLOCK(pll_lock),
        .O_LOCK(lock),
        .ICPSEL(icpsel),
        .LPFRES(lpfres)
    );
    defparam u_pll_init_HDMI.CLK_PERIOD = 20;
    defparam u_pll_init_HDMI.MULTI_FAC = 16;


endmodule
